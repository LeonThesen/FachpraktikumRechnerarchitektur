--
-- VHDL Architecture RISCV_Processor_lib.dbpu.behav
--
-- Created:
--          by - st161569.st161569 (pc043)
--          at - 17:26:57 05/29/24
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--
ARCHITECTURE behav OF dbpu IS
BEGIN
END ARCHITECTURE behav;

